`timescale 1ns / 1ps

module top #(
    parameter  IMEM_DEPTH = 4,       
    parameter  REGF_WIDTH = 16,     
    parameter  ALU_WIDTH = 16,       
    parameter  PROG_VALUE = 3

    );
    
      
  
  
  
endmodule


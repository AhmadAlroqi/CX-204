`timescale 1ns / 1ps


module alu  #(parameter int ALU_WIDTH = 16 ) 
(

    );
endmodule
